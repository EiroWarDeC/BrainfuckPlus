module main

fn main() {
	// 定义变量：操作的列表
	mut list_ptr := u32(0)
	mut list := []u8{len: 3000, cap: 3000, init: 0}
	// 定义变量：操作的代码字符串
	mut code_ptr := int(0)

	// 开始输出
	println('这是BrainfuckPlus的命令行运行程序，该程序使用V语言开发')
}